`timescale 1 ns / 1 ps

module AESL_deadlock_detector (
    input reset,
    input clock);

    wire [0:0] proc_dep_vld_vec_0;
    reg [0:0] proc_dep_vld_vec_0_reg;
    wire [0:0] in_chan_dep_vld_vec_0;
    wire [3:0] in_chan_dep_data_vec_0;
    wire [0:0] token_in_vec_0;
    wire [0:0] out_chan_dep_vld_vec_0;
    wire [3:0] out_chan_dep_data_0;
    wire [0:0] token_out_vec_0;
    wire dl_detect_out_0;
    wire dep_chan_vld_1_0;
    wire [3:0] dep_chan_data_1_0;
    wire token_1_0;
    wire [1:0] proc_dep_vld_vec_1;
    reg [1:0] proc_dep_vld_vec_1_reg;
    wire [1:0] in_chan_dep_vld_vec_1;
    wire [7:0] in_chan_dep_data_vec_1;
    wire [1:0] token_in_vec_1;
    wire [1:0] out_chan_dep_vld_vec_1;
    wire [3:0] out_chan_dep_data_1;
    wire [1:0] token_out_vec_1;
    wire dl_detect_out_1;
    wire dep_chan_vld_0_1;
    wire [3:0] dep_chan_data_0_1;
    wire token_0_1;
    wire dep_chan_vld_2_1;
    wire [3:0] dep_chan_data_2_1;
    wire token_2_1;
    wire [1:0] proc_dep_vld_vec_2;
    reg [1:0] proc_dep_vld_vec_2_reg;
    wire [1:0] in_chan_dep_vld_vec_2;
    wire [7:0] in_chan_dep_data_vec_2;
    wire [1:0] token_in_vec_2;
    wire [1:0] out_chan_dep_vld_vec_2;
    wire [3:0] out_chan_dep_data_2;
    wire [1:0] token_out_vec_2;
    wire dl_detect_out_2;
    wire dep_chan_vld_1_2;
    wire [3:0] dep_chan_data_1_2;
    wire token_1_2;
    wire dep_chan_vld_3_2;
    wire [3:0] dep_chan_data_3_2;
    wire token_3_2;
    wire [0:0] proc_dep_vld_vec_3;
    reg [0:0] proc_dep_vld_vec_3_reg;
    wire [0:0] in_chan_dep_vld_vec_3;
    wire [3:0] in_chan_dep_data_vec_3;
    wire [0:0] token_in_vec_3;
    wire [0:0] out_chan_dep_vld_vec_3;
    wire [3:0] out_chan_dep_data_3;
    wire [0:0] token_out_vec_3;
    wire dl_detect_out_3;
    wire dep_chan_vld_2_3;
    wire [3:0] dep_chan_data_2_3;
    wire token_2_3;
    wire [3:0] dl_in_vec;
    wire dl_detect_out;
    wire [3:0] origin;
    wire token_clear;

    reg ap_done_reg_0;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_0 <= 'b0;
        end
        else begin
            ap_done_reg_0 <= AESL_inst_MUSIC_top.inputdatamover_U0.ap_done;
        end
    end

    reg ap_done_reg_1;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_1 <= 'b0;
        end
        else begin
            ap_done_reg_1 <= AESL_inst_MUSIC_top.AutoCorrelation_U0.ap_done;
        end
    end

    reg ap_done_reg_2;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_2 <= 'b0;
        end
        else begin
            ap_done_reg_2 <= AESL_inst_MUSIC_top.qr_givens_U0.ap_done;
        end
    end

    reg ap_done_reg_3;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_3 <= 'b0;
        end
        else begin
            ap_done_reg_3 <= AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_done;
        end
    end

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_MUSIC_top$inputdatamover_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_MUSIC_top$inputdatamover_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_MUSIC_top$inputdatamover_U0$ap_idle <= AESL_inst_MUSIC_top.inputdatamover_U0.ap_idle;
        end
    end
    // Process: AESL_inst_MUSIC_top.inputdatamover_U0
    AESL_deadlock_detect_unit #(4, 0, 1, 1) AESL_deadlock_detect_unit_0 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_0),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_0),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_0),
        .token_in_vec(token_in_vec_0),
        .dl_detect_in(dl_detect_out),
        .origin(origin[0]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_0),
        .out_chan_dep_data(out_chan_dep_data_0),
        .token_out_vec(token_out_vec_0),
        .dl_detect_out(dl_in_vec[0]));

    assign proc_dep_vld_vec_0[0] = dl_detect_out ? proc_dep_vld_vec_0_reg[0] : (~AESL_inst_MUSIC_top.inMAT_re_U.i_full_n & AESL_inst_MUSIC_top.inputdatamover_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_MUSIC_top.inMAT_re_U.t_read | ~AESL_inst_MUSIC_top.inMAT_im_U.i_full_n & AESL_inst_MUSIC_top.inputdatamover_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_MUSIC_top.inMAT_im_U.t_read);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_0_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_0_reg <= proc_dep_vld_vec_0;
        end
    end
    assign in_chan_dep_vld_vec_0[0] = dep_chan_vld_1_0;
    assign in_chan_dep_data_vec_0[3 : 0] = dep_chan_data_1_0;
    assign token_in_vec_0[0] = token_1_0;
    assign dep_chan_vld_0_1 = out_chan_dep_vld_vec_0[0];
    assign dep_chan_data_0_1 = out_chan_dep_data_0;
    assign token_0_1 = token_out_vec_0[0];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_MUSIC_top$AutoCorrelation_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_MUSIC_top$AutoCorrelation_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_MUSIC_top$AutoCorrelation_U0$ap_idle <= AESL_inst_MUSIC_top.AutoCorrelation_U0.ap_idle;
        end
    end
    // Process: AESL_inst_MUSIC_top.AutoCorrelation_U0
    AESL_deadlock_detect_unit #(4, 1, 2, 2) AESL_deadlock_detect_unit_1 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_1),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_1),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_1),
        .token_in_vec(token_in_vec_1),
        .dl_detect_in(dl_detect_out),
        .origin(origin[1]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_1),
        .out_chan_dep_data(out_chan_dep_data_1),
        .token_out_vec(token_out_vec_1),
        .dl_detect_out(dl_in_vec[1]));

    assign proc_dep_vld_vec_1[0] = dl_detect_out ? proc_dep_vld_vec_1_reg[0] : (~AESL_inst_MUSIC_top.inMAT_re_U.t_empty_n & (AESL_inst_MUSIC_top.AutoCorrelation_U0.ap_ready | AESL_inst_MUSIC_top.AutoCorrelation_U0.ap_idle) & ~AESL_inst_MUSIC_top.inMAT_re_U.i_write | ~AESL_inst_MUSIC_top.inMAT_im_U.t_empty_n & (AESL_inst_MUSIC_top.AutoCorrelation_U0.ap_ready | AESL_inst_MUSIC_top.AutoCorrelation_U0.ap_idle) & ~AESL_inst_MUSIC_top.inMAT_im_U.i_write);
    assign proc_dep_vld_vec_1[1] = dl_detect_out ? proc_dep_vld_vec_1_reg[1] : (~AESL_inst_MUSIC_top.matrix1_re_U.i_full_n & AESL_inst_MUSIC_top.AutoCorrelation_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_MUSIC_top.matrix1_re_U.t_read | ~AESL_inst_MUSIC_top.matrix1_im_U.i_full_n & AESL_inst_MUSIC_top.AutoCorrelation_U0.ap_done & deadlock_detector.ap_done_reg_1 & ~AESL_inst_MUSIC_top.matrix1_im_U.t_read);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_1_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_1_reg <= proc_dep_vld_vec_1;
        end
    end
    assign in_chan_dep_vld_vec_1[0] = dep_chan_vld_0_1;
    assign in_chan_dep_data_vec_1[3 : 0] = dep_chan_data_0_1;
    assign token_in_vec_1[0] = token_0_1;
    assign in_chan_dep_vld_vec_1[1] = dep_chan_vld_2_1;
    assign in_chan_dep_data_vec_1[7 : 4] = dep_chan_data_2_1;
    assign token_in_vec_1[1] = token_2_1;
    assign dep_chan_vld_1_0 = out_chan_dep_vld_vec_1[0];
    assign dep_chan_data_1_0 = out_chan_dep_data_1;
    assign token_1_0 = token_out_vec_1[0];
    assign dep_chan_vld_1_2 = out_chan_dep_vld_vec_1[1];
    assign dep_chan_data_1_2 = out_chan_dep_data_1;
    assign token_1_2 = token_out_vec_1[1];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_MUSIC_top$qr_givens_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_MUSIC_top$qr_givens_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_MUSIC_top$qr_givens_U0$ap_idle <= AESL_inst_MUSIC_top.qr_givens_U0.ap_idle;
        end
    end
    // Process: AESL_inst_MUSIC_top.qr_givens_U0
    AESL_deadlock_detect_unit #(4, 2, 2, 2) AESL_deadlock_detect_unit_2 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_2),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_2),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_2),
        .token_in_vec(token_in_vec_2),
        .dl_detect_in(dl_detect_out),
        .origin(origin[2]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_2),
        .out_chan_dep_data(out_chan_dep_data_2),
        .token_out_vec(token_out_vec_2),
        .dl_detect_out(dl_in_vec[2]));

    assign proc_dep_vld_vec_2[0] = dl_detect_out ? proc_dep_vld_vec_2_reg[0] : (~AESL_inst_MUSIC_top.matrix1_re_U.t_empty_n & (AESL_inst_MUSIC_top.qr_givens_U0.ap_ready | AESL_inst_MUSIC_top.qr_givens_U0.ap_idle) & ~AESL_inst_MUSIC_top.matrix1_re_U.i_write | ~AESL_inst_MUSIC_top.matrix1_im_U.t_empty_n & (AESL_inst_MUSIC_top.qr_givens_U0.ap_ready | AESL_inst_MUSIC_top.qr_givens_U0.ap_idle) & ~AESL_inst_MUSIC_top.matrix1_im_U.i_write);
    assign proc_dep_vld_vec_2[1] = dl_detect_out ? proc_dep_vld_vec_2_reg[1] : (~AESL_inst_MUSIC_top.noiseSS_0_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_0_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_1_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_1_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_2_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_2_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_3_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_3_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_4_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_4_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_5_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_5_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_6_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_6_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_7_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_7_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_8_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_8_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_9_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_9_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_10_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_10_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_11_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_11_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_12_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_12_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_13_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_13_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_14_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_14_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_15_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_15_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_16_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_16_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_17_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_17_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_18_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_18_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_19_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_19_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_20_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_20_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_21_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_21_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_22_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_22_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_23_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_23_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_24_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_24_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_25_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_25_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_26_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_26_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_27_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_27_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_28_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_28_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_29_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_29_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_30_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_30_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_31_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_31_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_32_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_32_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_33_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_33_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_34_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_34_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_35_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_35_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_36_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_36_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_37_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_37_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_38_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_38_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_39_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_39_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_40_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_40_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_41_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_41_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_42_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_42_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_43_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_43_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_44_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_44_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_45_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_45_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_46_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_46_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_47_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_47_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_48_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_48_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_49_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_49_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_50_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_50_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_51_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_51_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_52_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_52_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_53_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_53_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_54_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_54_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_55_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_55_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_56_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_56_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_57_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_57_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_58_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_58_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_59_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_59_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_60_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_60_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_61_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_61_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_62_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_62_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_63_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_63_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_64_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_64_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_65_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_65_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_66_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_66_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_67_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_67_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_68_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_68_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_69_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_69_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_70_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_70_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_71_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_71_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_72_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_72_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_73_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_73_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_74_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_74_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_75_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_75_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_76_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_76_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_77_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_77_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_78_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_78_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_79_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_79_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_80_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_80_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_81_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_81_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_82_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_82_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_83_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_83_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_84_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_84_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_85_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_85_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_86_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_86_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_87_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_87_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_88_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_88_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_89_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_89_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_90_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_90_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_91_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_91_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_92_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_92_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_93_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_93_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_94_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_94_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_95_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_95_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_96_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_96_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_97_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_97_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_98_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_98_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_99_re_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_99_re_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_0_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_0_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_1_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_1_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_2_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_2_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_3_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_3_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_4_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_4_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_5_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_5_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_6_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_6_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_7_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_7_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_8_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_8_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_9_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_9_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_10_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_10_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_11_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_11_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_12_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_12_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_13_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_13_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_14_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_14_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_15_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_15_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_16_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_16_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_17_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_17_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_18_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_18_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_19_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_19_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_20_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_20_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_21_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_21_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_22_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_22_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_23_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_23_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_24_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_24_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_25_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_25_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_26_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_26_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_27_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_27_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_28_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_28_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_29_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_29_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_30_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_30_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_31_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_31_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_32_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_32_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_33_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_33_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_34_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_34_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_35_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_35_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_36_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_36_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_37_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_37_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_38_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_38_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_39_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_39_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_40_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_40_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_41_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_41_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_42_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_42_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_43_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_43_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_44_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_44_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_45_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_45_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_46_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_46_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_47_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_47_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_48_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_48_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_49_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_49_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_50_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_50_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_51_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_51_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_52_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_52_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_53_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_53_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_54_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_54_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_55_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_55_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_56_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_56_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_57_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_57_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_58_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_58_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_59_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_59_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_60_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_60_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_61_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_61_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_62_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_62_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_63_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_63_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_64_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_64_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_65_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_65_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_66_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_66_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_67_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_67_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_68_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_68_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_69_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_69_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_70_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_70_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_71_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_71_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_72_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_72_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_73_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_73_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_74_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_74_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_75_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_75_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_76_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_76_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_77_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_77_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_78_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_78_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_79_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_79_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_80_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_80_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_81_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_81_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_82_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_82_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_83_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_83_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_84_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_84_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_85_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_85_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_86_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_86_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_87_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_87_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_88_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_88_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_89_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_89_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_90_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_90_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_91_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_91_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_92_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_92_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_93_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_93_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_94_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_94_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_95_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_95_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_96_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_96_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_97_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_97_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_98_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_98_im_U.t_read | ~AESL_inst_MUSIC_top.noiseSS_99_im_U.i_full_n & AESL_inst_MUSIC_top.qr_givens_U0.ap_done & deadlock_detector.ap_done_reg_2 & ~AESL_inst_MUSIC_top.noiseSS_99_im_U.t_read);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_2_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_2_reg <= proc_dep_vld_vec_2;
        end
    end
    assign in_chan_dep_vld_vec_2[0] = dep_chan_vld_1_2;
    assign in_chan_dep_data_vec_2[3 : 0] = dep_chan_data_1_2;
    assign token_in_vec_2[0] = token_1_2;
    assign in_chan_dep_vld_vec_2[1] = dep_chan_vld_3_2;
    assign in_chan_dep_data_vec_2[7 : 4] = dep_chan_data_3_2;
    assign token_in_vec_2[1] = token_3_2;
    assign dep_chan_vld_2_1 = out_chan_dep_vld_vec_2[0];
    assign dep_chan_data_2_1 = out_chan_dep_data_2;
    assign token_2_1 = token_out_vec_2[0];
    assign dep_chan_vld_2_3 = out_chan_dep_vld_vec_2[1];
    assign dep_chan_data_2_3 = out_chan_dep_data_2;
    assign token_2_3 = token_out_vec_2[1];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_MUSIC_top$MSG_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_MUSIC_top$MSG_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_MUSIC_top$MSG_U0$ap_idle <= AESL_inst_MUSIC_top.MSG_U0.ap_idle;
        end
    end
    // Process: AESL_inst_MUSIC_top.MSG_U0
    AESL_deadlock_detect_unit #(4, 3, 1, 1) AESL_deadlock_detect_unit_3 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_3),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_3),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_3),
        .token_in_vec(token_in_vec_3),
        .dl_detect_in(dl_detect_out),
        .origin(origin[3]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_3),
        .out_chan_dep_data(out_chan_dep_data_3),
        .token_out_vec(token_out_vec_3),
        .dl_detect_out(dl_in_vec[3]));

    assign proc_dep_vld_vec_3[0] = dl_detect_out ? proc_dep_vld_vec_3_reg[0] : (~AESL_inst_MUSIC_top.noiseSS_0_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_0_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_1_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_1_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_2_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_2_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_3_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_3_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_4_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_4_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_5_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_5_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_6_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_6_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_7_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_7_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_8_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_8_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_9_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_9_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_10_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_10_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_11_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_11_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_12_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_12_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_13_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_13_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_14_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_14_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_15_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_15_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_16_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_16_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_17_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_17_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_18_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_18_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_19_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_19_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_20_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_20_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_21_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_21_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_22_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_22_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_23_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_23_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_24_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_24_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_25_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_25_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_26_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_26_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_27_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_27_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_28_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_28_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_29_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_29_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_30_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_30_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_31_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_31_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_32_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_32_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_33_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_33_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_34_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_34_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_35_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_35_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_36_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_36_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_37_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_37_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_38_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_38_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_39_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_39_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_40_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_40_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_41_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_41_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_42_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_42_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_43_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_43_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_44_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_44_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_45_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_45_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_46_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_46_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_47_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_47_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_48_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_48_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_49_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_49_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_50_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_50_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_51_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_51_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_52_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_52_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_53_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_53_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_54_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_54_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_55_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_55_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_56_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_56_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_57_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_57_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_58_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_58_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_59_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_59_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_60_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_60_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_61_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_61_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_62_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_62_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_63_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_63_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_64_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_64_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_65_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_65_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_66_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_66_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_67_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_67_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_68_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_68_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_69_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_69_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_70_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_70_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_71_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_71_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_72_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_72_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_73_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_73_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_74_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_74_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_75_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_75_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_76_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_76_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_77_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_77_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_78_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_78_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_79_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_79_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_80_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_80_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_81_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_81_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_82_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_82_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_83_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_83_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_84_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_84_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_85_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_85_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_86_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_86_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_87_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_87_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_88_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_88_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_89_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_89_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_90_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_90_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_91_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_91_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_92_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_92_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_93_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_93_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_94_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_94_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_95_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_95_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_96_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_96_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_97_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_97_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_98_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_98_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_99_re_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_99_re_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_0_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_0_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_1_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_1_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_2_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_2_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_3_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_3_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_4_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_4_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_5_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_5_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_6_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_6_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_7_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_7_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_8_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_8_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_9_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_9_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_10_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_10_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_11_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_11_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_12_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_12_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_13_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_13_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_14_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_14_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_15_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_15_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_16_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_16_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_17_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_17_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_18_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_18_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_19_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_19_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_20_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_20_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_21_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_21_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_22_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_22_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_23_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_23_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_24_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_24_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_25_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_25_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_26_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_26_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_27_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_27_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_28_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_28_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_29_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_29_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_30_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_30_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_31_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_31_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_32_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_32_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_33_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_33_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_34_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_34_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_35_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_35_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_36_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_36_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_37_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_37_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_38_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_38_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_39_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_39_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_40_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_40_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_41_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_41_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_42_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_42_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_43_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_43_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_44_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_44_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_45_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_45_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_46_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_46_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_47_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_47_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_48_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_48_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_49_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_49_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_50_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_50_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_51_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_51_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_52_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_52_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_53_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_53_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_54_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_54_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_55_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_55_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_56_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_56_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_57_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_57_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_58_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_58_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_59_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_59_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_60_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_60_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_61_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_61_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_62_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_62_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_63_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_63_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_64_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_64_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_65_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_65_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_66_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_66_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_67_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_67_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_68_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_68_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_69_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_69_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_70_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_70_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_71_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_71_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_72_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_72_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_73_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_73_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_74_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_74_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_75_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_75_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_76_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_76_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_77_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_77_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_78_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_78_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_79_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_79_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_80_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_80_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_81_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_81_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_82_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_82_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_83_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_83_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_84_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_84_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_85_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_85_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_86_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_86_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_87_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_87_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_88_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_88_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_89_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_89_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_90_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_90_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_91_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_91_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_92_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_92_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_93_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_93_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_94_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_94_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_95_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_95_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_96_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_96_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_97_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_97_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_98_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_98_im_U.i_write | ~AESL_inst_MUSIC_top.noiseSS_99_im_U.t_empty_n & (AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_ready | AESL_inst_MUSIC_top.MSG_U0.grp_matmul2_fu_1721.ap_idle) & ~AESL_inst_MUSIC_top.noiseSS_99_im_U.i_write);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_3_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_3_reg <= proc_dep_vld_vec_3;
        end
    end
    assign in_chan_dep_vld_vec_3[0] = dep_chan_vld_2_3;
    assign in_chan_dep_data_vec_3[3 : 0] = dep_chan_data_2_3;
    assign token_in_vec_3[0] = token_2_3;
    assign dep_chan_vld_3_2 = out_chan_dep_vld_vec_3[0];
    assign dep_chan_data_3_2 = out_chan_dep_data_3;
    assign token_3_2 = token_out_vec_3[0];


    AESL_deadlock_report_unit #(4) AESL_deadlock_report_unit_inst (
        .reset(reset),
        .clock(clock),
        .dl_in_vec(dl_in_vec),
        .dl_detect_out(dl_detect_out),
        .origin(origin),
        .token_clear(token_clear));

endmodule
